module dm74ls85(
    input wire [7:4] a,
    input wire [7:4] b,
    output wire aeb, // a == b
    output wire agb, // a > b
    output wire alb  // a < b
);


endmodule